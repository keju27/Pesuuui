
// Write code for modules you need here

module alu (input wire [1:0] op, input wire [15:0] i0, i1,
    output wire [15:0] o, output wire cout);

// Declare wires here

// Instantiate modules here

endmodule
